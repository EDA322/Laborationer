LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY EDA322_processor IS	Port (	       externalIn 	  : IN  std_logic_vector (7 DOWNTO 0);  -- “extIn” in Figure 1	       CLK 		  : IN  std_logic;	       master_load_enable : IN  std_logic;	       ARESETN 	   	  : IN  std_logic;	       pc2seg 	 	  : OUT std_logic_vector (7 DOWNTO 0);  -- PC	       instr2seg 	  : OUT std_logic_vector (11 DOWNTO 0); -- Instruction register	       Addr2seg   	  : OUT std_logic_vector (7 DOWNTO 0);  -- Address register	       dMemOut2seg 	  : OUT std_logic_vector (7 DOWNTO 0);  -- Data memory output	       aluOut2seg  	  : OUT std_logic_vector (7 DOWNTO 0);  -- ALU output	       acc2seg 	   	  : OUT std_logic_vector (7 DOWNTO 0);  -- Accumulator	       flag2seg    	  : OUT std_logic_vector (3 DOWNTO 0);  -- Flags	       busOut2seg  	  : OUT std_logic_vector (7 DOWNTO 0);  -- Value on the bus	       disp2seg   	  : OUT std_logic_vector(7 DOWNTO 0);   -- Display register	       errSig2seg  	  : OUT std_logic;                      -- Bus Error signal	       ovf	   	  : OUT std_logic;                      -- Overflow	       zero 	   	  : OUT std_logic);                     -- ZeroEND EDA322_processor;