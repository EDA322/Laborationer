LIBRARY ieee;USE ieee.std_logic_1164.all;USE ieee.numeric_std.all;

PACKAGE procComponents ISCOMPONENT procController    Port ( master_load_enable: in STD_LOGIC;	   opcode : in  STD_LOGIC_VECTOR (3 downto 0);	   neq : in STD_LOGIC;	   eq : in STD_LOGIC; 	   CLK : in STD_LOGIC;           ARESETN : in STD_LOGIC;	   pcSel : out  STD_LOGIC;	   pcLd : out  STD_LOGIC;	   instrLd : out  STD_LOGIC;	   addrMd : out  STD_LOGIC;           dmWr : out  STD_LOGIC;	   dataLd : out  STD_LOGIC;	   flagLd : out  STD_LOGIC;	   accSel : out  STD_LOGIC;	   accLd : out  STD_LOGIC;	   im2bus : out  STD_LOGIC;	   dmRd : out  STD_LOGIC;	   acc2bus : out  STD_LOGIC;	   ext2bus : out  STD_LOGIC;	   dispLd: out STD_LOGIC;	   aluMd : out STD_LOGIC_VECTOR(1 downto 0)
	);END COMPONENT;COMPONENT procBus    PORT ( INSTRUCTION : IN  std_logic_vector (7 DOWNTO 0);           DATA	       : IN  std_logic_vector (7 DOWNTO 0);           ACC 	       : IN  std_logic_vector (7 DOWNTO 0);           EXTDATA     : IN  std_logic_vector (7 DOWNTO 0);           OUTPUT      : OUT std_logic_vector (7 DOWNTO 0);           ERR         : OUT std_logic;           instrSEL    : IN  std_logic;           dataSEL     : IN  std_logic;           accSEL      : IN  std_logic;           extdataSEL  : IN  std_logic
	);END COMPONENT;COMPONENT alu_wRCA	PORT( ALU_inA, ALU_inB : in STD_LOGIC_VECTOR(7 downto 0);	      Operation : in STD_LOGIC_VECTOR(1 downto 0);	      ALU_out : out STD_LOGIC_VECTOR(7 downto 0);	      Carry, NotEq, Eq, isOutZero : out STD_LOGIC
	);END COMPONENT;COMPONENT alu_wCLA	PORT( ALU_inA, ALU_inB : in STD_LOGIC_VECTOR(7 downto 0);	      Operation : in STD_LOGIC_VECTOR(1 downto 0);	      ALU_out : out STD_LOGIC_VECTOR(7 downto 0);	      Carry, NotEq, Eq, isOutZero : out STD_LOGIC
	);END COMPONENT;COMPONENT mux2to1	GENERIC ( width: integer:=8);	PORT ( w1 : in STD_LOGIC_VECTOR(width-1 downto 0);	       w2 : in STD_LOGIC_VECTOR(width-1 downto 0);		       f : out STD_LOGIC_VECTOR(width-1 downto 0);		       sel : in STD_LOGIC
	);END COMPONENT;COMPONENT mem_array	GENERIC ( DATA_WIDTH : integer := 12;		  ADDR_WIDTH : integer := 8;		  INIT_FILE  : string  := "inst_mem.mif");	PORT ( ADDR    : IN STD_LOGIC_VECTOR (ADDR_WIDTH-1 DOWNTO 0);	       DATA_IN : IN STD_LOGIC_VECTOR (DATA_WIDTH-1 DOWNTO 0);	       CLK     : IN STD_LOGIC;	       WE      : IN STD_LOGIC;	       OUTPUT  : OUT STD_LOGIC_VECTOR (DATA_WIDTH-1 DOWNTO 0)
	);END COMPONENT;COMPONENT reg	GENERIC( width: integer := 8 );	PORT( CLK 	 : IN std_logic;	      ARESETN	 : IN std_logic;	      loadEnable : IN std_logic;	      input      : IN std_logic_vector(width-1 DOWNTO 0);	      res        : OUT std_logic_vector(width-1 DOWNTO 0)	);END COMPONENT;END procComponents;