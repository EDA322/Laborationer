library ieee;use ieee.std_logic_1164.all;use ieee.numeric_std.all;

package procComponents IScomponent procController  port (  master_load_enable  : in std_logic;          opcode              : in std_logic_vector (3 downto 0);          neq                 : in std_logic;          eq                  : in std_logic;          CLK                 : in std_logic;          ARESETN             : in std_logic;          pcSel               : out std_logic;          pcLd                : out std_logic;          instrLd             : out std_logic;          addrMd              : out std_logic;          dmWr                : out std_logic;          dataLd              : out std_logic;          flagLd              : out std_logic;          accSel              : out std_logic;          accLd               : out std_logic;          im2bus              : out std_logic;          dmRd                : out std_logic;          acc2bus             : out std_logic;          ext2bus             : out std_logic;          dispLd              : out std_logic;          aluMd               : out std_logic_vector(1 downto 0) );
end component;component procBus  port (  INSTRUCTION         : in  std_logic_vector (7 downto 0);          DATA	              : in  std_logic_vector (7 downto 0);          ACC 	              : in  std_logic_vector (7 downto 0);          EXTDATA             : in  std_logic_vector (7 downto 0);          OUTPUT              : out std_logic_vector (7 downto 0);          ERR                 : out std_logic;          instrSEL            : in  std_logic;          dataSEL             : in  std_logic;          accSEL              : in  std_logic;          extdataSEL          : in  std_logic );
end component;component alu_wRCA  port (  ALU_inA, ALU_inB      : in std_logic_vector(7 downto 0);	        Operation             : in std_logic_vector(1 downto 0);	        ALU_out               : out std_logic_vector(7 downto 0);	        Carry, NotEq, Eq      : out std_logic;
          isOutZero             : out std_logic );
end component;component alu_wCLA	port (  ALU_inA, ALU_inB      : in std_logic_vector(7 downto 0);	        Operation             : in std_logic_vector(1 downto 0);	        ALU_out               : out std_logic_vector(7 downto 0);	        Carry, NotEq, Eq      : out std_logic;
          isOutZero             : out std_logic );
end component;component mux2to1	generic (  width: integer:=8);	port (  w1                    : in std_logic_vector(width-1 downto 0);	        w2                    : in std_logic_vector(width-1 downto 0);          f                     : out std_logic_vector(width-1 downto 0);          sel                   : in std_logic  );
end component;component mem_array	generic (  DATA_WIDTH : integer := 12;		         ADDR_WIDTH : integer := 8;		         INIT_FILE  : string  := "inst_mem.mif" );	port (  ADDR                  : in std_logic_vector(ADDR_WIDTH-1 downto 0);	        DATA_IN               : in std_logic_vector(DATA_WIDTH-1 downto 0);	        CLK                   : in std_logic;	        WE                    : in std_logic;	        OUTPUT                : out std_logic_vector(DATA_WIDTH-1 downto 0) );
end component;component reg	generic (  width: integer := 8 );	port (  CLK 	                : in std_logic;	        ARESETN	              : in std_logic;	        loadEnable            : in std_logic;  	      input                 : in std_logic_vector(width-1 downto 0);  	      res                   : out std_logic_vector(width-1 downto 0) );end component;end procComponents;